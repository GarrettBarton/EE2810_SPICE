Hor_2_39
*E	+	-	val
*VIN 1	0	DC 0.5V
XP	6	5	1	POT PARAMS: R=10K SET={SET}
X1	0	2	5	6	3	UA741
*+INPUT	-INPUT +VCC -VEE OUTPUT CONNECTIONS FOR UA741
VCC 5	0	15V
VEE	6	0	-15V
R1	1	2	1500
R2	2	3	1000
**************************
*(TOP, BOTTOM, TAP)
.SUBCKT POT 6 5 1 PARAMS: VALUE=10K SET=0.5
RT 6 1 {VALUE*(1-SET)+.001}
RB 1 5 {VALUE*SET+.001}
.ENDS
**************************
*.DC VIN -15 +15 .5V
.TRAN 0.1ms 1s
.PARAM SET=.5
.STEP PARAM(SET) 0, 1, .2
.LIB NOM.LIB
.PROBE V(3)
.END